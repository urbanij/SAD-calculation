---------------------------------------------
-- Title       : tb_SAD_wrapper
-- Project     : Final project: SAD Calculation
---------------------------------------------
-- File        : tb_SAD_wrapper.vhd
-- Language    : VHDL
-- Author(s)   : Francesco Urbani
-- Company     : 
-- Created     : Sun May 27 20:53:15 CEST 2018
---------------------------------------------
-- Description : Autogenerated test bench for SAD.vhd
---------------------------------------------
-- Update      :
---------------------------------------------

-- THIS TEST BENCH IS AUTOGENERATED FROM SAD_model.py
-- WARNING! All changes made in this file might be lost!



-- INPUTS:
-- N  = 8 bits
-- px = 16

-- SAD_bits_min := min num bits to correctly represent SAD
-- SAD_bits_min = ceil( log2( (2**N-1) * px**2 )) = 
--              = ceil( log2( 255 * 256 )) = 
--              = 16


-- PA = 
--     [249 129 148 110  82   6 186 195 125   0  31 100 235 231  55 222]
--     [ 83 125 123  32 143  17  95 216  77 143 159 252 137 228  81 124]
--     [219 232   2  63  40  69 155   7  71  80 190 236 191 188   1  54]
--     [ 72 137  68 186 100 106 175 208 238 123  56 244 216  91 108 232]
--     [ 24  83  83  26  87 212  86  67  60 231   7  27 242 106  34 249]
--     [129 120 136 221 118 232 238   0 200  88 172 216   7 168 149 240]
--     [  6  52 208 244 121   9  40 118 174  34  67  26 138 187  27 208]
--     [188  28 216 111 189 136  43  99 116 162  24 149  59 124 107 194]
--     [111  40   8 145 139  45 249 188 198 168  36   3 244 244 104 162]
--     [144  79 205  78 119 186  85 203 113 221   0  11 194 193 143 116]
--     [193  60  20  66 173 128 156 126 213  17 238 172 239 110 155 210]
--     [114 230 251  56  63  88 112   5   8 124 122 229  72 134  79 160]
--     [154 135 113  61  42  53  26  58 220  15  31 229 191 149 127 141]
--     [ 87  70 139 223  67 168  32  91 135  83  42 154  24 151 156 147]
--     [133 201 181  71  76 228  43 247  61  60 242 168 237  94  65 228]
--     [  7 174  41  19 131 200 235 233 152 174 223  85  12 201  79 158]
-- PB = 
--     [ 12  67  91 250 182 208 137 248   1 213 123 225 176  66   5 253]
--     [142 132 172  36 179 168 108  78  61 247 134  58 220  26  33 227]
--     [245  31 245 126 248 171 178 123  96 195 115   1 187 236 114  73]
--     [ 62  49 252 134   2 250 106 107 127  74  30 156  88 240 134  47]
--     [132  92 253 108  35  71 242 255 198  19  98  68 252  46  48 111]
--     [236 116  17 177  40 165  57 237  40 170 176  43 106  32 121 232]
--     [219  42  57  37   3 133  16 251  48  56 255 211  32 155 185  58]
--     [ 23  16 232 110  60 126 117 134 176  69  94 149 193 192 107 224]
--     [251  69  35 199  42  20  80 217 175 203 168   0 215 200  83  63]
--     [103  23 178 158  68 233 115 219   6  16 251 122 139 209 120  79]
--     [227 175 119  11 220 209  92 143 109  26  13  48  39  15 184 123]
--     [132  51 131 226  71  10 212 159 212  46  98 209  67  78 222 122]
--     [ 65  19  29  12  61  76  95  56 107 180 191 232 116 189  18 129]
--     [199 131  76 161 147   1 122 133  49  15 177 196  33 242 149  94]
--     [  0  41 178  98 196 253 239  91 180 162 197 110  12 209  58  84]
--     [ 44 173 123  60 108  16 144  63 124 197  78  68 103  60 189 121]

-- OUTPUT:
-- DIFF = 
--     [237  62  57 140 100 202  49  53 124 213  92 125  59 165  50  31]
--     [ 59   7  49   4  36 151  13 138  16 104  25 194  83 202  48 103]
--     [ 26 201 243  63 208 102  23 116  25 115  75 235   4  48 113  19]
--     [ 10  88 184  52  98 144  69 101 111  49  26  88 128 149  26 185]
--     [108   9 170  82  52 141 156 188 138 212  91  41  10  60  14 138]
--     [107   4 119  44  78  67 181 237 160  82   4 173  99 136  28   8]
--     [213  10 151 207 118 124  24 133 126  22 188 185 106  32 158 150]
--     [165  12  16   1 129  10  74  35  60  93  70   0 134  68   0  30]
--     [140  29  27  54  97  25 169  29  23  35 132   3  29  44  21  99]
--     [ 41  56  27  80  51  47  30  16 107 205 251 111  55  16  23  37]
--     [ 34 115  99  55  47  81  64  17 104   9 225 124 200  95  29  87]
--     [ 18 179 120 170   8  78 100 154 204  78  24  20   5  56 143  38]
--     [ 89 116  84  49  19  23  69   2 113 165 160   3  75  40 109  12]
--     [112  61  63  62  80 167  90  42  86  68 135  42   9  91   7  53]
--     [133 160   3  27 120  25 196 156 119 102  45  58 225 115   7 144]
--     [ 37   1  82  41  23 184  91 170  28  23 145  17  91 141 110  37]

-- SAD_value = sum(SAD) = 22137 = "0101011001111001"



library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;


entity tb_SAD_wrapper is
end entity tb_SAD_wrapper; -- tb_SAD_wrapper


architecture struct of tb_SAD_wrapper is
	
	component SAD is
		generic(
			Npixel     : positive ;      -- total # of pixels of the image
			
			Nbit       : positive ;        -- # of bits needed to represent the value of each pixel
			SAD_bits   : positive  	-- # of bits needed to represent the output
		);
		port(
			CLK        : in  std_logic;
			RST        : in  std_logic;
			EN         : in  std_logic;
			PA         : in  std_logic_vector(Nbit-1  downto 0);
			PB         : in  std_logic_vector(Nbit-1  downto 0);
			
			SAD        : out std_logic_vector(SAD_bits-1 downto 0); 
			DATA_VALID : out std_logic
		);
	end component SAD;


	constant Npixel  : positive := 256;
	constant Nbit    : positive := 8;
	constant Mbit    : positive := 16;
	constant clk_per : time     := 5 ns;

	signal clk       : std_logic := '0';
	signal reset     : std_logic ;
	signal enable    : std_logic ;
	signal PA        : std_logic_vector(Nbit-1 downto 0) := "00000000";
	signal PB        : std_logic_vector(Nbit-1 downto 0) := "XXXXXXXX";

	signal sad : std_logic_vector(M-1 downto 0);
	signal DATA_VALID: std_logic;


	signal testing   : Boolean   := True;




begin
	clk <= not clk after clk_per/2 when testing;-- ELSE '0';


	sad_i: SAD_wrapper
		generic map(Npixel, Nbit, Mbit)
		port map(clk, reset, enable, PA, PB, sad, DATA_VALID);


	drive_p: process
	  	begin
			
			
			PA <= "01000001";
			PB <= "11000011";
			wait until rising_edge(clk);

			PA <= "01110001";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "01101100";
			PB <= "01010000";
			wait until rising_edge(clk);

			PA <= "00011101";
			PB <= "01011000";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "10100001";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "00111011";
			wait until rising_edge(clk);

			PA <= "01001110";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "11001101";
			PB <= "01101001";
			wait until rising_edge(clk);

			PA <= "10011001";
			PB <= "11100111";
			wait until rising_edge(clk);

			PA <= "00000000";
			PB <= "00000000";
			wait until rising_edge(clk);

-----------------------


			PA <= "11111001";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "01000011";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "01010010";
			PB <= "10110110";
			wait until rising_edge(clk);

			PA <= "00000110";
			PB <= "11010000";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "10001001";
			wait until rising_edge(clk);

			PA <= "11000011";
			PB <= "11111000";
			wait until rising_edge(clk);

			PA <= "01111101";
			PB <= "00000001";
			wait until rising_edge(clk);

			PA <= "00000000";
			PB <= "11010101";
			wait until rising_edge(clk);

			PA <= "00011111";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "01100100";
			PB <= "11100001";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "10110000";
			wait until rising_edge(clk);

			PA <= "11100111";
			PB <= "01000010";
			wait until rising_edge(clk);

			PA <= "00110111";
			PB <= "00000101";
			wait until rising_edge(clk);

			PA <= "11011110";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "01111101";
			PB <= "10000100";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "10101100";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "10001111";
			PB <= "10110011";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "01011111";
			PB <= "01101100";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "01001101";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "10001111";
			PB <= "11110111";
			wait until rising_edge(clk);

			PA <= "10011111";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "11111100";
			PB <= "00111010";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "11100100";
			PB <= "00011010";
			wait until rising_edge(clk);

			PA <= "01010001";
			PB <= "00100001";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "00011111";
			wait until rising_edge(clk);

			PA <= "00000010";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "00111111";
			PB <= "01111110";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "11111000";
			wait until rising_edge(clk);

			PA <= "01000101";
			PB <= "10101011";
			wait until rising_edge(clk);

			PA <= "10011011";
			PB <= "10110010";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "01100000";
			wait until rising_edge(clk);

			PA <= "01010000";
			PB <= "11000011";
			wait until rising_edge(clk);

			PA <= "10111110";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "00000001";
			wait until rising_edge(clk);

			PA <= "10111111";
			PB <= "10111011";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "11101100";
			wait until rising_edge(clk);

			PA <= "00000001";
			PB <= "01110010";
			wait until rising_edge(clk);

			PA <= "00110110";
			PB <= "01001001";
			wait until rising_edge(clk);

			PA <= "01001000";
			PB <= "00111110";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "01000100";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "01100100";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "01101010";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "01101010";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "01101011";
			wait until rising_edge(clk);

			PA <= "11101110";
			PB <= "01111111";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "01001010";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "11110100";
			PB <= "10011100";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "01011000";
			wait until rising_edge(clk);

			PA <= "01011011";
			PB <= "11110000";
			wait until rising_edge(clk);

			PA <= "01101100";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "00101111";
			wait until rising_edge(clk);

			PA <= "00011000";
			PB <= "10000100";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "01011100";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "00011010";
			PB <= "01101100";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "00100011";
			wait until rising_edge(clk);

			PA <= "11010100";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "01010110";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "01000011";
			PB <= "11111111";
			wait until rising_edge(clk);

			PA <= "00111100";
			PB <= "11000110";
			wait until rising_edge(clk);

			PA <= "11100111";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01100010";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "11110010";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "01101010";
			PB <= "00101110";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "00110000";
			wait until rising_edge(clk);

			PA <= "11111001";
			PB <= "01101111";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "11101100";
			wait until rising_edge(clk);

			PA <= "01111000";
			PB <= "01110100";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "00010001";
			wait until rising_edge(clk);

			PA <= "11011101";
			PB <= "10110001";
			wait until rising_edge(clk);

			PA <= "01110110";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "10100101";
			wait until rising_edge(clk);

			PA <= "11101110";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "00000000";
			PB <= "11101101";
			wait until rising_edge(clk);

			PA <= "11001000";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "10101010";
			wait until rising_edge(clk);

			PA <= "10101100";
			PB <= "10110000";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01101010";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "10010101";
			PB <= "01111001";
			wait until rising_edge(clk);

			PA <= "11110000";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "00000110";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "11110100";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "01111001";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "00001001";
			PB <= "10000101";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "01110110";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "10101110";
			PB <= "00110000";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "00111000";
			wait until rising_edge(clk);

			PA <= "01000011";
			PB <= "11111111";
			wait until rising_edge(clk);

			PA <= "00011010";
			PB <= "11010011";
			wait until rising_edge(clk);

			PA <= "10001010";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "10111011";
			PB <= "10011011";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "10111001";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "00111010";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "00010111";
			wait until rising_edge(clk);

			PA <= "00011100";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "10111101";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "01111110";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "01110101";
			wait until rising_edge(clk);

			PA <= "01100011";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "01110100";
			PB <= "10110000";
			wait until rising_edge(clk);

			PA <= "10100010";
			PB <= "01000101";
			wait until rising_edge(clk);

			PA <= "00011000";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "10010101";
			PB <= "10010101";
			wait until rising_edge(clk);

			PA <= "00111011";
			PB <= "11000001";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "11000000";
			wait until rising_edge(clk);

			PA <= "01101011";
			PB <= "01101011";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "01000101";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "00100011";
			wait until rising_edge(clk);

			PA <= "10010001";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "10001011";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "00101101";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "11111001";
			PB <= "01010000";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "11011001";
			wait until rising_edge(clk);

			PA <= "11000110";
			PB <= "10101111";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "11001011";
			wait until rising_edge(clk);

			PA <= "00100100";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "00000011";
			PB <= "00000000";
			wait until rising_edge(clk);

			PA <= "11110100";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "11110100";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "01101000";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "10100010";
			PB <= "00111111";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "01100111";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "00010111";
			wait until rising_edge(clk);

			PA <= "11001101";
			PB <= "10110010";
			wait until rising_edge(clk);

			PA <= "01001110";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "01110111";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "11101001";
			wait until rising_edge(clk);

			PA <= "01010101";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "01110001";
			PB <= "00000110";
			wait until rising_edge(clk);

			PA <= "11011101";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "00000000";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "00001011";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "10001011";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "10001111";
			PB <= "01111000";
			wait until rising_edge(clk);

			PA <= "01110100";
			PB <= "01001111";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "00111100";
			PB <= "10101111";
			wait until rising_edge(clk);

			PA <= "00010100";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "01000010";
			PB <= "00001011";
			wait until rising_edge(clk);

			PA <= "10101101";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "01011100";
			wait until rising_edge(clk);

			PA <= "01111110";
			PB <= "10001111";
			wait until rising_edge(clk);

			PA <= "11010101";
			PB <= "01101101";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "00011010";
			wait until rising_edge(clk);

			PA <= "11101110";
			PB <= "00001101";
			wait until rising_edge(clk);

			PA <= "10101100";
			PB <= "00110000";
			wait until rising_edge(clk);

			PA <= "11101111";
			PB <= "00100111";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "10011011";
			PB <= "10111000";
			wait until rising_edge(clk);

			PA <= "11010010";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "10000100";
			wait until rising_edge(clk);

			PA <= "11100110";
			PB <= "00110011";
			wait until rising_edge(clk);

			PA <= "11111011";
			PB <= "10000011";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "11100010";
			wait until rising_edge(clk);

			PA <= "00111111";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "01110000";
			PB <= "11010100";
			wait until rising_edge(clk);

			PA <= "00000101";
			PB <= "10011111";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "11010100";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "00101110";
			wait until rising_edge(clk);

			PA <= "01111010";
			PB <= "01100010";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "01001000";
			PB <= "01000011";
			wait until rising_edge(clk);

			PA <= "10000110";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "11011110";
			wait until rising_edge(clk);

			PA <= "10100000";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "10000111";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "01110001";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "00111101";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "00110101";
			PB <= "01001100";
			wait until rising_edge(clk);

			PA <= "00011010";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "00111010";
			PB <= "00111000";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "01101011";
			wait until rising_edge(clk);

			PA <= "00001111";
			PB <= "10110100";
			wait until rising_edge(clk);

			PA <= "00011111";
			PB <= "10111111";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "10111111";
			PB <= "01110100";
			wait until rising_edge(clk);

			PA <= "10010101";
			PB <= "10111101";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "00010010";
			wait until rising_edge(clk);

			PA <= "10001101";
			PB <= "10000001";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "10000011";
			wait until rising_edge(clk);

			PA <= "10001011";
			PB <= "01001100";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "10100001";
			wait until rising_edge(clk);

			PA <= "01000011";
			PB <= "10010011";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "00000001";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "01011011";
			PB <= "10000101";
			wait until rising_edge(clk);

			PA <= "10000111";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "10110001";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "11000100";
			wait until rising_edge(clk);

			PA <= "00011000";
			PB <= "00100001";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "10010101";
			wait until rising_edge(clk);

			PA <= "10010011";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "10000101";
			PB <= "00000000";
			wait until rising_edge(clk);

			PA <= "11001001";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "10110101";
			PB <= "10110010";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "01100010";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "11000100";
			wait until rising_edge(clk);

			PA <= "11100100";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "00111101";
			PB <= "10110100";
			wait until rising_edge(clk);

			PA <= "00111100";
			PB <= "10100010";
			wait until rising_edge(clk);

			PA <= "11110010";
			PB <= "11000101";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "11101101";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "00111010";
			wait until rising_edge(clk);

			PA <= "11100100";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "10101110";
			PB <= "10101101";
			wait until rising_edge(clk);

			PA <= "00101001";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "00010011";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "10000011";
			PB <= "01101100";
			wait until rising_edge(clk);

			PA <= "11001000";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "10010000";
			wait until rising_edge(clk);

			PA <= "11101001";
			PB <= "00111111";
			wait until rising_edge(clk);

			PA <= "10011000";
			PB <= "01111100";
			wait until rising_edge(clk);

			PA <= "10101110";
			PB <= "11000101";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "01010101";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "01100111";
			wait until rising_edge(clk);

			PA <= "11001001";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "10111101";
			wait until rising_edge(clk);

			PA <= "10011110";
			PB <= "01111001";
			wait until rising_edge(clk);


------------------------------------------


			PA <= "01011001";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "10011000";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "11010001";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "10001110";
			PB <= "00110110";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "10011001";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "01100111";
			PB <= "00110101";
			wait until rising_edge(clk);

			PA <= "01100001";
			PB <= "10000011";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "00110010";
			PB <= "00000111";
			wait until rising_edge(clk);

			PA <= "11011010";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "11101010";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "01111101";
			wait until rising_edge(clk);

			PA <= "11010010";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "11101101";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "00000010";
			PB <= "10000101";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "11001111";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "00111111";
			wait until rising_edge(clk);

			PA <= "00101100";
			PB <= "01100110";
			wait until rising_edge(clk);

			PA <= "01101000";
			PB <= "11110000";
			wait until rising_edge(clk);

			PA <= "11010100";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "10100111";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "01111001";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "01110101";
			PB <= "10001100";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "00101110";
			PB <= "01011010";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "00001010";
			PB <= "00011001";
			wait until rising_edge(clk);

			PA <= "01110011";
			PB <= "11000001";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "00010101";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "01010000";
			PB <= "00000110";
			wait until rising_edge(clk);

			PA <= "10110111";
			PB <= "00001001";
			wait until rising_edge(clk);

			PA <= "01110110";
			PB <= "00100111";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "01000000";
			wait until rising_edge(clk);

			PA <= "01111010";
			PB <= "11001010";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "10110111";
			wait until rising_edge(clk);

			PA <= "00010010";
			PB <= "10010011";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "11101110";
			wait until rising_edge(clk);

			PA <= "11010010";
			PB <= "10111110";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "01111111";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "10101101";
			wait until rising_edge(clk);

			PA <= "11000101";
			PB <= "01101011";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "01001000";
			PB <= "01010101";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "11101100";
			wait until rising_edge(clk);

			PA <= "00110101";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "00000101";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "11001001";
			wait until rising_edge(clk);

			PA <= "11111110";
			PB <= "10000001";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "01011010";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "01001001";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "00110010";
			wait until rising_edge(clk);

			PA <= "00100110";
			PB <= "10011101";
			wait until rising_edge(clk);

			PA <= "00001011";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "11011101";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "01100111";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "10111110";
			PB <= "11110100";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "11010110";
			PB <= "10000111";
			wait until rising_edge(clk);

			PA <= "00000010";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "10110110";
			PB <= "10000000";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "01000101";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "10110000";
			wait until rising_edge(clk);

			PA <= "01101101";
			PB <= "11001010";
			wait until rising_edge(clk);

			PA <= "01010001";
			PB <= "11011110";
			wait until rising_edge(clk);

			PA <= "00111101";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "11101101";
			wait until rising_edge(clk);

			PA <= "10111001";
			PB <= "01111000";
			wait until rising_edge(clk);

			PA <= "00010111";
			PB <= "11101110";
			wait until rising_edge(clk);

			PA <= "00001110";
			PB <= "00011100";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "01011100";
			wait until rising_edge(clk);

			PA <= "01010001";
			PB <= "10110100";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "10110011";
			PB <= "00001110";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "10000100";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "10011111";
			PB <= "01000110";
			wait until rising_edge(clk);

			PA <= "10110100";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "11101111";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "01100110";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "10011111";
			PB <= "11100110";
			wait until rising_edge(clk);

			PA <= "00001110";
			PB <= "10010010";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "10011111";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "11001111";
			wait until rising_edge(clk);

			PA <= "11110011";
			PB <= "10011010";
			wait until rising_edge(clk);

			PA <= "00110011";
			PB <= "10111101";
			wait until rising_edge(clk);

			PA <= "10111111";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "00111110";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "11101101";
			PB <= "00110011";
			wait until rising_edge(clk);

			PA <= "11001100";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "01100010";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "01110111";
			PB <= "10010000";
			wait until rising_edge(clk);

			PA <= "10011011";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "10110010";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "11100010";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "00110101";
			PB <= "11000010";
			wait until rising_edge(clk);

			PA <= "11111111";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "00001010";
			PB <= "00111111";
			wait until rising_edge(clk);

			PA <= "10001111";
			PB <= "11110111";
			wait until rising_edge(clk);

			PA <= "00100100";
			PB <= "10100100";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "00010000";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "11101010";
			wait until rising_edge(clk);

			PA <= "10010110";
			PB <= "10111110";
			wait until rising_edge(clk);

			PA <= "10000110";
			PB <= "01110101";
			wait until rising_edge(clk);

			PA <= "10110110";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "00011111";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "10111011";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "00000101";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "00100001";
			wait until rising_edge(clk);

			PA <= "01110110";
			PB <= "10000011";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "01101010";
			wait until rising_edge(clk);

			PA <= "10111001";
			PB <= "01111001";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "11000000";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "00111010";
			PB <= "00000101";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "11111000";
			wait until rising_edge(clk);

			PA <= "10111000";
			PB <= "00011000";
			wait until rising_edge(clk);

			PA <= "11001001";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "10110110";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "11000010";
			wait until rising_edge(clk);

			PA <= "10111001";
			PB <= "11100100";
			wait until rising_edge(clk);

			PA <= "11111011";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "01110001";
			PB <= "00010010";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "11110110";
			wait until rising_edge(clk);

			PA <= "10100001";
			PB <= "10111000";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "11011000";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "10110110";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "11110011";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "01100011";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "00111111";
			PB <= "00101110";
			wait until rising_edge(clk);

			PA <= "10010101";
			PB <= "11011010";
			wait until rising_edge(clk);

			PA <= "11010100";
			PB <= "10001001";
			wait until rising_edge(clk);

			PA <= "10001011";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "10010001";
			PB <= "00011111";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "11000010";
			wait until rising_edge(clk);

			PA <= "00110000";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "10011111";
			PB <= "11110000";
			wait until rising_edge(clk);

			PA <= "01100000";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "11110001";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "01010010";
			wait until rising_edge(clk);

			PA <= "01010010";
			PB <= "11000010";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "01010111";
			wait until rising_edge(clk);

			PA <= "00001101";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "10001011";
			wait until rising_edge(clk);

			PA <= "10110111";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "01100111";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "01100000";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "01000000";
			PB <= "11110110";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "11010110";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "01111001";
			wait until rising_edge(clk);

			PA <= "10101110";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "01100101";
			PB <= "11100100";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "11111111";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "01110100";
			wait until rising_edge(clk);

			PA <= "01101011";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "01011101";
			PB <= "00110111";
			wait until rising_edge(clk);

			PA <= "10101100";
			PB <= "10001101";
			wait until rising_edge(clk);

			PA <= "01110100";
			PB <= "11101010";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "01100101";
			wait until rising_edge(clk);

			PA <= "01110111";
			PB <= "01001100";
			wait until rising_edge(clk);

			PA <= "11010001";
			PB <= "01001100";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "11100100";
			wait until rising_edge(clk);

			PA <= "00110101";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "00110000";
			PB <= "10111001";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "10100000";
			PB <= "00001001";
			wait until rising_edge(clk);

			PA <= "00100110";
			PB <= "11010101";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "10101100";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "01001111";
			wait until rising_edge(clk);

			PA <= "01110101";
			PB <= "10111011";
			wait until rising_edge(clk);

			PA <= "11101010";
			PB <= "10111001";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "00100011";
			wait until rising_edge(clk);

			PA <= "01000000";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "11100110";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "00101111";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "10111001";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "00000110";
			PB <= "11010011";
			wait until rising_edge(clk);

			PA <= "11011010";
			PB <= "11001010";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "00011010";
			wait until rising_edge(clk);

			PA <= "01010110";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "00011001";
			wait until rising_edge(clk);

			PA <= "10000010";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "11010011";
			PB <= "11001101";
			wait until rising_edge(clk);

			PA <= "01111110";
			PB <= "01011100";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "11111111";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "01010001";
			wait until rising_edge(clk);

			PA <= "01100111";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "10110101";
			PB <= "01011010";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "00000111";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "11000100";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "00000100";
			PB <= "10101100";
			wait until rising_edge(clk);

			PA <= "11111000";
			PB <= "01111111";
			wait until rising_edge(clk);

			PA <= "01111110";
			PB <= "00100010";
			wait until rising_edge(clk);

			PA <= "01001010";
			PB <= "10101100";
			wait until rising_edge(clk);

			PA <= "10111110";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "00010101";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "01011001";
			PB <= "01101111";
			wait until rising_edge(clk);

			PA <= "11000110";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "11000100";
			wait until rising_edge(clk);

			PA <= "00110101";
			PB <= "01010001";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "11011110";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "10010111";
			wait until rising_edge(clk);

			PA <= "10101101";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "10110100";
			PB <= "10111100";
			wait until rising_edge(clk);

			PA <= "11010111";
			PB <= "01111101";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "11001011";
			wait until rising_edge(clk);

			PA <= "10000101";
			PB <= "10001010";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "11001110";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "01100101";
			wait until rising_edge(clk);

			PA <= "00111111";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "00100110";
			PB <= "10000111";
			wait until rising_edge(clk);

			PA <= "00000001";
			PB <= "11000101";
			wait until rising_edge(clk);

			PA <= "11001111";
			PB <= "01111001";
			wait until rising_edge(clk);

			PA <= "10111011";
			PB <= "01000011";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "00001110";
			PB <= "01101101";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "10011010";
			wait until rising_edge(clk);

			PA <= "10100100";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "00100001";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "10101001";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "00001101";
			wait until rising_edge(clk);

			PA <= "11111111";
			PB <= "00010011";
			wait until rising_edge(clk);


------------------------------------------


			PA <= "00001110";
			PB <= "11111001";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "01001111";
			wait until rising_edge(clk);

			PA <= "00010011";
			PB <= "11011101";
			wait until rising_edge(clk);

			PA <= "01110100";
			PB <= "01001001";
			wait until rising_edge(clk);

			PA <= "11101010";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "10100000";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "01010010";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "00011100";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "11010110";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "01000010";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "11100000";
			PB <= "11010110";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "11000011";
			PB <= "10010101";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "00110100";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "01111110";
			wait until rising_edge(clk);

			PA <= "00001110";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "11110101";
			PB <= "11001010";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "00101110";
			wait until rising_edge(clk);

			PA <= "10001110";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "01011100";
			PB <= "10010111";
			wait until rising_edge(clk);

			PA <= "01000011";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "10010110";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "00010001";
			wait until rising_edge(clk);

			PA <= "00011001";
			PB <= "01001011";
			wait until rising_edge(clk);

			PA <= "11110011";
			PB <= "11000011";
			wait until rising_edge(clk);

			PA <= "10000010";
			PB <= "11101010";
			wait until rising_edge(clk);

			PA <= "00111011";
			PB <= "10100111";
			wait until rising_edge(clk);

			PA <= "10111000";
			PB <= "10110011";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "01110010";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "01100000";
			PB <= "10011010";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "00110110";
			wait until rising_edge(clk);

			PA <= "01011101";
			PB <= "11011101";
			wait until rising_edge(clk);

			PA <= "00010011";
			PB <= "10001000";
			wait until rising_edge(clk);

			PA <= "01111010";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "01100000";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "10011100";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "00001001";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "10001100";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "00011101";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "10111000";
			PB <= "00010001";
			wait until rising_edge(clk);

			PA <= "10010010";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "11111110";
			PB <= "11111111";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "11000101";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "01000101";
			wait until rising_edge(clk);

			PA <= "11110101";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "11010001";
			PB <= "10011001";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "10111110";
			wait until rising_edge(clk);

			PA <= "00001101";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "10101111";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "00011100";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "11001101";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "01011010";
			wait until rising_edge(clk);

			PA <= "00011010";
			PB <= "00110000";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "00010010";
			wait until rising_edge(clk);

			PA <= "11111010";
			PB <= "10111100";
			wait until rising_edge(clk);

			PA <= "10100110";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "11001110";
			PB <= "10011100";
			wait until rising_edge(clk);

			PA <= "11001100";
			PB <= "10111111";
			wait until rising_edge(clk);

			PA <= "10000110";
			PB <= "00110111";
			wait until rising_edge(clk);

			PA <= "10110111";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "01110000";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "10100100";
			PB <= "11110011";
			wait until rising_edge(clk);

			PA <= "10100101";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "11101010";
			wait until rising_edge(clk);

			PA <= "00101001";
			PB <= "11010000";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "00011000";
			wait until rising_edge(clk);

			PA <= "11001111";
			PB <= "11010010";
			wait until rising_edge(clk);

			PA <= "00011001";
			PB <= "11111110";
			wait until rising_edge(clk);

			PA <= "00001110";
			PB <= "00010010";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "00011010";
			PB <= "01110110";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "11000101";
			wait until rising_edge(clk);

			PA <= "10110110";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "10001010";
			wait until rising_edge(clk);

			PA <= "00111100";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "10011001";
			PB <= "01100110";
			wait until rising_edge(clk);

			PA <= "10010001";
			PB <= "10001101";
			wait until rising_edge(clk);

			PA <= "10111011";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "00011001";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "10010100";
			wait until rising_edge(clk);

			PA <= "00101100";
			PB <= "10101010";
			wait until rising_edge(clk);

			PA <= "01100010";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "10010010";
			wait until rising_edge(clk);

			PA <= "01011101";
			PB <= "01000000";
			wait until rising_edge(clk);

			PA <= "01111000";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "01000100";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "00111011";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "00000001";
			PB <= "01110100";
			wait until rising_edge(clk);

			PA <= "00011000";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "01010101";
			PB <= "11101110";
			wait until rising_edge(clk);

			PA <= "11001000";
			PB <= "00000111";
			wait until rising_edge(clk);

			PA <= "01011001";
			PB <= "10000001";
			wait until rising_edge(clk);

			PA <= "01110011";
			PB <= "10111001";
			wait until rising_edge(clk);

			PA <= "11110011";
			PB <= "00000001";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "00001011";
			wait until rising_edge(clk);

			PA <= "10110011";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "11010001";
			PB <= "00010010";
			wait until rising_edge(clk);

			PA <= "11110000";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "11110101";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "10110001";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "01010010";
			PB <= "10110111";
			wait until rising_edge(clk);

			PA <= "00001011";
			PB <= "11000011";
			wait until rising_edge(clk);

			PA <= "10000011";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "00010000";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "10010101";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "01100110";
			PB <= "01101100";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "01001001";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "01011101";
			wait until rising_edge(clk);

			PA <= "00101111";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "11110011";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "01001101";
			wait until rising_edge(clk);

			PA <= "10110010";
			PB <= "11111000";
			wait until rising_edge(clk);

			PA <= "01100100";
			PB <= "10001011";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "10001101";
			PB <= "10001111";
			wait until rising_edge(clk);

			PA <= "10001110";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "11110011";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "11101101";
			wait until rising_edge(clk);

			PA <= "11011110";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "00100100";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "00000101";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "00000110";
			PB <= "11110100";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "01111001";
			PB <= "01010101";
			wait until rising_edge(clk);

			PA <= "01110110";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "00100111";
			PB <= "11010100";
			wait until rising_edge(clk);

			PA <= "01100010";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "11110110";
			PB <= "00001011";
			wait until rising_edge(clk);

			PA <= "10100100";
			PB <= "11110011";
			wait until rising_edge(clk);

			PA <= "10001111";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "11001110";
			wait until rising_edge(clk);

			PA <= "01110011";
			PB <= "00110110";
			wait until rising_edge(clk);

			PA <= "01101011";
			PB <= "10100111";
			wait until rising_edge(clk);

			PA <= "01001011";
			PB <= "00001101";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "00001000";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "01100010";
			wait until rising_edge(clk);

			PA <= "11100000";
			PB <= "01111000";
			wait until rising_edge(clk);

			PA <= "10010110";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "10010100";
			wait until rising_edge(clk);

			PA <= "00011110";
			PB <= "01010101";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "10110000";
			wait until rising_edge(clk);

			PA <= "01110000";
			PB <= "11100100";
			wait until rising_edge(clk);

			PA <= "01011011";
			PB <= "10101100";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "10000001";
			wait until rising_edge(clk);

			PA <= "00110010";
			PB <= "00011000";
			wait until rising_edge(clk);

			PA <= "01110011";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "11001101";
			PB <= "11001101";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "00000100";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "01001010";
			PB <= "01010111";
			wait until rising_edge(clk);

			PA <= "11111001";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "01100001";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "11011001";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "11100010";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "10000010";
			PB <= "11001010";
			wait until rising_edge(clk);

			PA <= "00011000";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "10001011";
			wait until rising_edge(clk);

			PA <= "01100101";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "01100010";
			wait until rising_edge(clk);

			PA <= "00010000";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "11111010";
			PB <= "01010000";
			wait until rising_edge(clk);

			PA <= "10010110";
			PB <= "10111110";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "00000100";
			wait until rising_edge(clk);

			PA <= "11000101";
			PB <= "00001011";
			wait until rising_edge(clk);

			PA <= "11001100";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "01000110";
			wait until rising_edge(clk);

			PA <= "00011100";
			PB <= "01010001";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "11110110";
			wait until rising_edge(clk);

			PA <= "00010011";
			PB <= "01100101";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "01101010";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "10011000";
			wait until rising_edge(clk);

			PA <= "11100000";
			PB <= "11010000";
			wait until rising_edge(clk);

			PA <= "10110100";
			PB <= "11000001";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "01101111";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "11100100";
			wait until rising_edge(clk);

			PA <= "11100011";
			PB <= "11010110";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "10000101";
			wait until rising_edge(clk);

			PA <= "00000011";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "01111000";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "01110000";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "10110101";
			wait until rising_edge(clk);

			PA <= "11100001";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "00011110";
			PB <= "10110001";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "10011101";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "11011000";
			wait until rising_edge(clk);

			PA <= "11100011";
			PB <= "11111110";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "10110010";
			PB <= "11110000";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "10011101";
			wait until rising_edge(clk);

			PA <= "11001000";
			PB <= "00111010";
			wait until rising_edge(clk);

			PA <= "01001011";
			PB <= "11101011";
			wait until rising_edge(clk);

			PA <= "01010101";
			PB <= "11100100";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "00000101";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "11000100";
			wait until rising_edge(clk);

			PA <= "01000010";
			PB <= "10110110";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "10101101";
			wait until rising_edge(clk);

			PA <= "11101111";
			PB <= "00011001";
			wait until rising_edge(clk);

			PA <= "10100101";
			PB <= "01100000";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "01101111";
			wait until rising_edge(clk);

			PA <= "11111000";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "11010011";
			wait until rising_edge(clk);

			PA <= "10101010";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "01001010";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "11001101";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "11011010";
			PB <= "00011000";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "10110101";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "10100010";
			wait until rising_edge(clk);

			PA <= "10001100";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "00000001";
			PB <= "00011010";
			wait until rising_edge(clk);

			PA <= "01111001";
			PB <= "00011010";
			wait until rising_edge(clk);

			PA <= "11100001";
			PB <= "01110010";
			wait until rising_edge(clk);

			PA <= "11110110";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "00001110";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "01101111";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "10101001";
			wait until rising_edge(clk);

			PA <= "01111110";
			PB <= "01001100";
			wait until rising_edge(clk);

			PA <= "11100110";
			PB <= "11000000";
			wait until rising_edge(clk);

			PA <= "01100110";
			PB <= "00010111";
			wait until rising_edge(clk);

			PA <= "00011010";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "00101111";
			PB <= "10111110";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "10101101";
			wait until rising_edge(clk);

			PA <= "01001010";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "00110111";
			PB <= "11101001";
			wait until rising_edge(clk);

			PA <= "11110010";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "11100111";
			PB <= "00100011";
			wait until rising_edge(clk);

			PA <= "00111010";
			PB <= "01011101";
			wait until rising_edge(clk);

			PA <= "01110101";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "01001101";
			PB <= "10000001";
			wait until rising_edge(clk);

			PA <= "11110010";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "10110100";
			wait until rising_edge(clk);

			PA <= "00010100";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "01000011";
			PB <= "11100001";
			wait until rising_edge(clk);

			PA <= "01010001";
			PB <= "00110111";
			wait until rising_edge(clk);

			PA <= "10001010";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "11001110";
			wait until rising_edge(clk);

			PA <= "11100011";
			PB <= "11000000";
			wait until rising_edge(clk);


------------------------------------------


			PA <= "10111000";
			PB <= "10111011";
			wait until rising_edge(clk);

			PA <= "10110101";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "01001001";
			PB <= "10010100";
			wait until rising_edge(clk);

			PA <= "01000111";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "11000000";
			PB <= "10101011";
			wait until rising_edge(clk);

			PA <= "10100000";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "00011111";
			PB <= "10100001";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "01001010";
			wait until rising_edge(clk);

			PA <= "11001110";
			PB <= "00010111";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "01011101";
			wait until rising_edge(clk);

			PA <= "11001101";
			PB <= "11101110";
			wait until rising_edge(clk);

			PA <= "00000011";
			PB <= "10100111";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "10010010";
			PB <= "10010010";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "10010011";
			PB <= "11010100";
			wait until rising_edge(clk);

			PA <= "11110000";
			PB <= "10110101";
			wait until rising_edge(clk);

			PA <= "00001010";
			PB <= "00010110";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "10111100";
			wait until rising_edge(clk);

			PA <= "00110111";
			PB <= "11001001";
			wait until rising_edge(clk);

			PA <= "00001011";
			PB <= "10110111";
			wait until rising_edge(clk);

			PA <= "00000100";
			PB <= "10110011";
			wait until rising_edge(clk);

			PA <= "01100000";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "01001001";
			wait until rising_edge(clk);

			PA <= "01000101";
			PB <= "00011001";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "10001011";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "01101000";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "11011101";
			PB <= "01100110";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "10010011";
			wait until rising_edge(clk);

			PA <= "11110110";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "00100001";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "11000001";
			wait until rising_edge(clk);

			PA <= "00011001";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "10111010";
			PB <= "10101000";
			wait until rising_edge(clk);

			PA <= "10111011";
			PB <= "01110000";
			wait until rising_edge(clk);

			PA <= "00110000";
			PB <= "11110110";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "01100001";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "00100101";
			wait until rising_edge(clk);

			PA <= "11010100";
			PB <= "01110001";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "11010011";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "11111001";
			PB <= "00110101";
			wait until rising_edge(clk);

			PA <= "00101101";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "01001001";
			PB <= "10110010";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "01101001";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "10100010";
			wait until rising_edge(clk);

			PA <= "00001010";
			PB <= "00111010";
			wait until rising_edge(clk);

			PA <= "00001101";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "11011111";
			wait until rising_edge(clk);

			PA <= "00110111";
			PB <= "11100001";
			wait until rising_edge(clk);

			PA <= "01001111";
			PB <= "01001011";
			wait until rising_edge(clk);

			PA <= "10001010";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "11101101";
			PB <= "10010010";
			wait until rising_edge(clk);

			PA <= "01101011";
			PB <= "10101110";
			wait until rising_edge(clk);

			PA <= "00100100";
			PB <= "00000110";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "11111001";
			PB <= "00100001";
			wait until rising_edge(clk);

			PA <= "00011100";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "10100110";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "00111001";
			PB <= "00110101";
			wait until rising_edge(clk);

			PA <= "10110100";
			PB <= "00111000";
			wait until rising_edge(clk);

			PA <= "00011111";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "01101001";
			wait until rising_edge(clk);

			PA <= "10010001";
			PB <= "10011101";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "01111000";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "10111111";
			wait until rising_edge(clk);

			PA <= "10001111";
			PB <= "11110110";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "11000010";
			wait until rising_edge(clk);

			PA <= "00101101";
			PB <= "00111011";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "01110000";
			wait until rising_edge(clk);

			PA <= "01100001";
			PB <= "00110110";
			wait until rising_edge(clk);

			PA <= "01010000";
			PB <= "10001000";
			wait until rising_edge(clk);

			PA <= "00000110";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "11100111";
			wait until rising_edge(clk);

			PA <= "10101011";
			PB <= "11111110";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "00011111";
			wait until rising_edge(clk);

			PA <= "10000010";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "00000100";
			PB <= "00011011";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "10010111";
			wait until rising_edge(clk);

			PA <= "10000100";
			PB <= "01000101";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "10001101";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "11100001";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "00111100";
			PB <= "11001111";
			wait until rising_edge(clk);

			PA <= "00001011";
			PB <= "01010111";
			wait until rising_edge(clk);

			PA <= "11111111";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "10001110";
			PB <= "10110110";
			wait until rising_edge(clk);

			PA <= "10100101";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "11000011";
			PB <= "00000001";
			wait until rising_edge(clk);

			PA <= "10111110";
			PB <= "11000110";
			wait until rising_edge(clk);

			PA <= "10011111";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "10100011";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "10101110";
			wait until rising_edge(clk);

			PA <= "10100111";
			PB <= "11000001";
			wait until rising_edge(clk);

			PA <= "11111001";
			PB <= "00110100";
			wait until rising_edge(clk);

			PA <= "00000010";
			PB <= "10001000";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "01011100";
			wait until rising_edge(clk);

			PA <= "11100000";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "10111001";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "01011000";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "00100011";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "00100010";
			wait until rising_edge(clk);

			PA <= "10011000";
			PB <= "11100010";
			wait until rising_edge(clk);

			PA <= "10100001";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "11000011";
			PB <= "01010101";
			wait until rising_edge(clk);

			PA <= "10111101";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "10010001";
			PB <= "10110001";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "10010100";
			wait until rising_edge(clk);

			PA <= "11100001";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "10110111";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "11100110";
			PB <= "00110011";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "10000000";
			wait until rising_edge(clk);

			PA <= "10010101";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "10110110";
			PB <= "01110101";
			wait until rising_edge(clk);

			PA <= "10010000";
			PB <= "01001011";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "01111101";
			wait until rising_edge(clk);

			PA <= "00010100";
			PB <= "10001001";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "01111110";
			wait until rising_edge(clk);

			PA <= "00101000";
			PB <= "00010110";
			wait until rising_edge(clk);

			PA <= "00101010";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "00111110";
			wait until rising_edge(clk);

			PA <= "10000110";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "11000000";
			PB <= "10001010";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "00001001";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "11010111";
			PB <= "11011001";
			wait until rising_edge(clk);

			PA <= "00110110";
			PB <= "00110011";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "01010100";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "00011011";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "01101101";
			PB <= "00011111";
			wait until rising_edge(clk);

			PA <= "00110001";
			PB <= "01111011";
			wait until rising_edge(clk);

			PA <= "00100100";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "00111001";
			PB <= "10000000";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "10001100";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "01000011";
			wait until rising_edge(clk);

			PA <= "10101110";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "10101000";
			PB <= "11000011";
			wait until rising_edge(clk);

			PA <= "00100011";
			PB <= "10001111";
			wait until rising_edge(clk);

			PA <= "10110111";
			PB <= "11110001";
			wait until rising_edge(clk);

			PA <= "00010010";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "11100001";
			PB <= "01110000";
			wait until rising_edge(clk);

			PA <= "10001101";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "00110101";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "00011101";
			PB <= "10001100";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "11101101";
			wait until rising_edge(clk);

			PA <= "00010100";
			PB <= "11111110";
			wait until rising_edge(clk);

			PA <= "00111100";
			PB <= "01111000";
			wait until rising_edge(clk);

			PA <= "01010000";
			PB <= "11100110";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "10101101";
			wait until rising_edge(clk);

			PA <= "01011100";
			PB <= "01001100";
			wait until rising_edge(clk);

			PA <= "01000010";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "00110111";
			PB <= "10001100";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "11010101";
			wait until rising_edge(clk);

			PA <= "01001110";
			PB <= "01110011";
			wait until rising_edge(clk);

			PA <= "11011000";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "10110110";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "01111001";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "11010000";
			wait until rising_edge(clk);

			PA <= "10001100";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "10011011";
			PB <= "10000100";
			wait until rising_edge(clk);

			PA <= "01111000";
			PB <= "01011001";
			wait until rising_edge(clk);

			PA <= "01110100";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "01111101";
			wait until rising_edge(clk);

			PA <= "10111101";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "11010110";
			PB <= "01001001";
			wait until rising_edge(clk);

			PA <= "01001000";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "00101101";
			wait until rising_edge(clk);

			PA <= "00010111";
			PB <= "00111011";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "10001010";
			PB <= "10001101";
			wait until rising_edge(clk);

			PA <= "11000101";
			PB <= "00111111";
			wait until rising_edge(clk);

			PA <= "00101101";
			PB <= "01010000";
			wait until rising_edge(clk);

			PA <= "10110100";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "11010010";
			PB <= "10010001";
			wait until rising_edge(clk);

			PA <= "01100111";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "10110001";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "10011011";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "00010011";
			PB <= "00010010";
			wait until rising_edge(clk);

			PA <= "10110010";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "11111000";
			PB <= "00001000";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "11101100";
			wait until rising_edge(clk);

			PA <= "10101100";
			PB <= "10100100";
			wait until rising_edge(clk);

			PA <= "01101100";
			PB <= "10110101";
			wait until rising_edge(clk);

			PA <= "01011011";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "01001101";
			PB <= "01011110";
			wait until rising_edge(clk);

			PA <= "00000110";
			PB <= "01001101";
			wait until rising_edge(clk);

			PA <= "11101001";
			PB <= "00111011";
			wait until rising_edge(clk);

			PA <= "01111010";
			PB <= "00101101";
			wait until rising_edge(clk);

			PA <= "01000011";
			PB <= "01100101";
			wait until rising_edge(clk);

			PA <= "01111101";
			PB <= "01000011";
			wait until rising_edge(clk);

			PA <= "11010100";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "10101011";
			wait until rising_edge(clk);

			PA <= "10110100";
			PB <= "01001101";
			wait until rising_edge(clk);

			PA <= "10110111";
			PB <= "11000000";
			wait until rising_edge(clk);

			PA <= "01000101";
			PB <= "01010101";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "00110100";
			wait until rising_edge(clk);

			PA <= "10111101";
			PB <= "10100100";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "10011111";
			wait until rising_edge(clk);

			PA <= "11011100";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "01001010";
			wait until rising_edge(clk);

			PA <= "10100101";
			PB <= "10000111";
			wait until rising_edge(clk);

			PA <= "00000010";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "00101110";
			wait until rising_edge(clk);

			PA <= "01010010";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "00011001";
			PB <= "00011001";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "10001000";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "01001011";
			wait until rising_edge(clk);

			PA <= "01000101";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "11101101";
			PB <= "11000011";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "00111001";
			wait until rising_edge(clk);

			PA <= "11010101";
			PB <= "10000010";
			wait until rising_edge(clk);

			PA <= "01000100";
			PB <= "01100101";
			wait until rising_edge(clk);

			PA <= "10100001";
			PB <= "10010011";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "00010001";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "01011010";
			PB <= "00001001";
			wait until rising_edge(clk);

			PA <= "11110110";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "10001001";
			wait until rising_edge(clk);

			PA <= "00110110";
			PB <= "01000110";
			wait until rising_edge(clk);

			PA <= "01001001";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "11100100";
			PB <= "10001001";
			wait until rising_edge(clk);

			PA <= "10110101";
			PB <= "11100110";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "00111000";
			wait until rising_edge(clk);

			PA <= "00011101";
			PB <= "10001011";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "11001100";
			PB <= "00011000";
			wait until rising_edge(clk);

			PA <= "01110111";
			PB <= "11111001";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "10000000";
			wait until rising_edge(clk);

			PA <= "01101001";
			PB <= "00011010";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "11011011";
			wait until rising_edge(clk);

			PA <= "10011110";
			PB <= "01110110";
			wait until rising_edge(clk);

			PA <= "10100000";
			PB <= "01111010";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "10001111";
			wait until rising_edge(clk);

			PA <= "11000100";
			PB <= "11101001";
			wait until rising_edge(clk);


------------------------------------------


			PA <= "00010100";
			PB <= "01000100";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "01000001";
			wait until rising_edge(clk);

			PA <= "10100011";
			PB <= "11101010";
			wait until rising_edge(clk);

			PA <= "00011111";
			PB <= "10101011";
			wait until rising_edge(clk);

			PA <= "10000100";
			PB <= "00011000";
			wait until rising_edge(clk);

			PA <= "11110111";
			PB <= "00000100";
			wait until rising_edge(clk);

			PA <= "01010101";
			PB <= "01100111";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "01001011";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "01011101";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "00001110";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "10101010";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "11011010";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "00110010";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "10010110";
			wait until rising_edge(clk);

			PA <= "10001101";
			PB <= "00000110";
			wait until rising_edge(clk);

			PA <= "10011001";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "00111000";
			wait until rising_edge(clk);

			PA <= "10000010";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "01111111";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "11101001";
			PB <= "01000110";
			wait until rising_edge(clk);

			PA <= "01000101";
			PB <= "10010100";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "01100100";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "11010001";
			wait until rising_edge(clk);

			PA <= "11011001";
			PB <= "10001101";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "11010111";
			wait until rising_edge(clk);

			PA <= "11101000";
			PB <= "11110000";
			wait until rising_edge(clk);

			PA <= "10100010";
			PB <= "11001101";
			wait until rising_edge(clk);

			PA <= "10101111";
			PB <= "10101110";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "00011101";
			PB <= "01000011";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "11100011";
			PB <= "11001111";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "10100110";
			PB <= "10010011";
			wait until rising_edge(clk);

			PA <= "00101100";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "11110000";
			wait until rising_edge(clk);

			PA <= "11101101";
			PB <= "11110001";
			wait until rising_edge(clk);

			PA <= "10001100";
			PB <= "11101110";
			wait until rising_edge(clk);

			PA <= "01100110";
			PB <= "10101010";
			wait until rising_edge(clk);

			PA <= "00011001";
			PB <= "00011111";
			wait until rising_edge(clk);

			PA <= "01111101";
			PB <= "10111100";
			wait until rising_edge(clk);

			PA <= "11010001";
			PB <= "01110000";
			wait until rising_edge(clk);

			PA <= "11001100";
			PB <= "11001110";
			wait until rising_edge(clk);

			PA <= "11101010";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "10100011";
			PB <= "10111000";
			wait until rising_edge(clk);

			PA <= "11111011";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "01110000";
			PB <= "10010010";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "01110100";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "00100111";
			wait until rising_edge(clk);

			PA <= "01100101";
			PB <= "00001110";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "00101111";
			PB <= "01011100";
			wait until rising_edge(clk);

			PA <= "10011000";
			PB <= "10011000";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "00100111";
			PB <= "00110000";
			wait until rising_edge(clk);

			PA <= "00101110";
			PB <= "00000100";
			wait until rising_edge(clk);

			PA <= "10011100";
			PB <= "11100111";
			wait until rising_edge(clk);

			PA <= "00101011";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "10010100";
			PB <= "01001101";
			wait until rising_edge(clk);

			PA <= "01001011";
			PB <= "11010011";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "10110100";
			wait until rising_edge(clk);

			PA <= "01000100";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "00011110";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "11011100";
			wait until rising_edge(clk);

			PA <= "11001100";
			PB <= "00010110";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "00110010";
			wait until rising_edge(clk);

			PA <= "11110001";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "10100000";
			wait until rising_edge(clk);

			PA <= "01001101";
			PB <= "10010101";
			wait until rising_edge(clk);

			PA <= "11001001";
			PB <= "10101111";
			wait until rising_edge(clk);

			PA <= "00111000";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "00010101";
			PB <= "00010011";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "00110010";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "11100111";
			wait until rising_edge(clk);

			PA <= "00111110";
			PB <= "11110001";
			wait until rising_edge(clk);

			PA <= "01001110";
			PB <= "00010110";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "10100101";
			PB <= "10100111";
			wait until rising_edge(clk);

			PA <= "10101010";
			PB <= "00100001";
			wait until rising_edge(clk);

			PA <= "00111110";
			PB <= "01110010";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "00000111";
			wait until rising_edge(clk);

			PA <= "10011000";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "10011000";
			PB <= "00001110";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "11011000";
			wait until rising_edge(clk);

			PA <= "00001011";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "10100111";
			PB <= "10101001";
			wait until rising_edge(clk);

			PA <= "01011010";
			PB <= "11110101";
			wait until rising_edge(clk);

			PA <= "00100011";
			PB <= "11100000";
			wait until rising_edge(clk);

			PA <= "10000100";
			PB <= "11101011";
			wait until rising_edge(clk);

			PA <= "10010111";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "01001001";
			PB <= "00101010";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "01001111";
			wait until rising_edge(clk);

			PA <= "00110110";
			PB <= "10110101";
			wait until rising_edge(clk);

			PA <= "10100011";
			PB <= "01110010";
			wait until rising_edge(clk);

			PA <= "11000011";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "10010011";
			PB <= "11000001";
			wait until rising_edge(clk);

			PA <= "10000010";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "01001011";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "10111100";
			PB <= "11110010";
			wait until rising_edge(clk);

			PA <= "00000100";
			PB <= "01110110";
			wait until rising_edge(clk);

			PA <= "10000001";
			PB <= "01010011";
			wait until rising_edge(clk);

			PA <= "01101011";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "01000010";
			PB <= "00000111";
			wait until rising_edge(clk);

			PA <= "11001111";
			PB <= "10011001";
			wait until rising_edge(clk);

			PA <= "00111111";
			PB <= "10011011";
			wait until rising_edge(clk);

			PA <= "01010100";
			PB <= "11111110";
			wait until rising_edge(clk);

			PA <= "01111110";
			PB <= "00100110";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "10111000";
			wait until rising_edge(clk);

			PA <= "00110100";
			PB <= "00010100";
			wait until rising_edge(clk);

			PA <= "11100100";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "10101110";
			PB <= "11100111";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "11101011";
			wait until rising_edge(clk);

			PA <= "11100100";
			PB <= "00001011";
			wait until rising_edge(clk);

			PA <= "11001001";
			PB <= "00110100";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "00001101";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "10011001";
			PB <= "01011010";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "01010000";
			wait until rising_edge(clk);

			PA <= "10011110";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "10000011";
			PB <= "10011011";
			wait until rising_edge(clk);

			PA <= "00010111";
			PB <= "00011011";
			wait until rising_edge(clk);

			PA <= "10011111";
			PB <= "01100110";
			wait until rising_edge(clk);

			PA <= "00011011";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "00000011";
			PB <= "11110001";
			wait until rising_edge(clk);

			PA <= "00101110";
			PB <= "10100100";
			wait until rising_edge(clk);

			PA <= "11111100";
			PB <= "00000010";
			wait until rising_edge(clk);

			PA <= "01001101";
			PB <= "11100101";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "11001011";
			wait until rising_edge(clk);

			PA <= "00101111";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "10111011";
			PB <= "11110100";
			wait until rising_edge(clk);

			PA <= "11100001";
			PB <= "00001101";
			wait until rising_edge(clk);

			PA <= "10100011";
			PB <= "00001000";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "10001101";
			wait until rising_edge(clk);

			PA <= "10100111";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "10001001";
			PB <= "00101000";
			wait until rising_edge(clk);

			PA <= "01110110";
			PB <= "11101111";
			wait until rising_edge(clk);

			PA <= "11011011";
			PB <= "11000000";
			wait until rising_edge(clk);

			PA <= "10001110";
			PB <= "10101011";
			wait until rising_edge(clk);

			PA <= "11111000";
			PB <= "00101001";
			wait until rising_edge(clk);

			PA <= "10101101";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "01101101";
			PB <= "10110010";
			wait until rising_edge(clk);

			PA <= "01011111";
			PB <= "10110100";
			wait until rising_edge(clk);

			PA <= "01001110";
			PB <= "01011010";
			wait until rising_edge(clk);

			PA <= "10110000";
			PB <= "10100101";
			wait until rising_edge(clk);

			PA <= "01101100";
			PB <= "10101110";
			wait until rising_edge(clk);

			PA <= "11100111";
			PB <= "10100011";
			wait until rising_edge(clk);

			PA <= "01100001";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "00000110";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "10101001";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "11111010";
			wait until rising_edge(clk);

			PA <= "00001010";
			PB <= "01101110";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "00010001";
			wait until rising_edge(clk);

			PA <= "00011000";
			PB <= "10001010";
			wait until rising_edge(clk);

			PA <= "00111011";
			PB <= "00111011";
			wait until rising_edge(clk);

			PA <= "11000001";
			PB <= "11000000";
			wait until rising_edge(clk);

			PA <= "10100101";
			PB <= "10111111";
			wait until rising_edge(clk);

			PA <= "11001000";
			PB <= "11010110";
			wait until rising_edge(clk);

			PA <= "10001011";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "01001100";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "01011011";
			wait until rising_edge(clk);

			PA <= "10000000";
			PB <= "00110001";
			wait until rising_edge(clk);

			PA <= "01001110";
			PB <= "00001100";
			wait until rising_edge(clk);

			PA <= "00110011";
			PB <= "01001111";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "11100000";
			PB <= "10110101";
			wait until rising_edge(clk);

			PA <= "01101101";
			PB <= "00111110";
			wait until rising_edge(clk);

			PA <= "00100010";
			PB <= "11011110";
			wait until rising_edge(clk);

			PA <= "11100010";
			PB <= "00100010";
			wait until rising_edge(clk);

			PA <= "11110101";
			PB <= "10111000";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "00001111";
			wait until rising_edge(clk);

			PA <= "01110010";
			PB <= "10000001";
			wait until rising_edge(clk);

			PA <= "01001011";
			PB <= "11111011";
			wait until rising_edge(clk);

			PA <= "00110000";
			PB <= "00101101";
			wait until rising_edge(clk);

			PA <= "01011101";
			PB <= "10100110";
			wait until rising_edge(clk);

			PA <= "11110001";
			PB <= "10100011";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "01110100";
			PB <= "11001100";
			wait until rising_edge(clk);

			PA <= "10000111";
			PB <= "11100011";
			wait until rising_edge(clk);

			PA <= "10111110";
			PB <= "10100101";
			wait until rising_edge(clk);

			PA <= "11001011";
			PB <= "01010101";
			wait until rising_edge(clk);

			PA <= "00101101";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "11110001";
			PB <= "01101100";
			wait until rising_edge(clk);

			PA <= "01111011";
			PB <= "01101111";
			wait until rising_edge(clk);

			PA <= "00010001";
			PB <= "10011001";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "10011101";
			PB <= "10000100";
			wait until rising_edge(clk);

			PA <= "11111110";
			PB <= "00001000";
			wait until rising_edge(clk);

			PA <= "00100001";
			PB <= "11000110";
			wait until rising_edge(clk);

			PA <= "00010110";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "01011101";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "11111101";
			PB <= "00011111";
			wait until rising_edge(clk);

			PA <= "01110001";
			PB <= "11100111";
			wait until rising_edge(clk);

			PA <= "01111100";
			PB <= "11111101";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "00100111";
			wait until rising_edge(clk);

			PA <= "01011111";
			PB <= "10111010";
			wait until rising_edge(clk);

			PA <= "01101111";
			PB <= "00111100";
			wait until rising_edge(clk);

			PA <= "01000001";
			PB <= "10111011";
			wait until rising_edge(clk);

			PA <= "11111011";
			PB <= "01111101";
			wait until rising_edge(clk);

			PA <= "10100110";
			PB <= "11101000";
			wait until rising_edge(clk);

			PA <= "01011110";
			PB <= "10011010";
			wait until rising_edge(clk);

			PA <= "11111011";
			PB <= "10110011";
			wait until rising_edge(clk);

			PA <= "10000110";
			PB <= "00000011";
			wait until rising_edge(clk);

			PA <= "11100101";
			PB <= "11110011";
			wait until rising_edge(clk);

			PA <= "00100100";
			PB <= "01001011";
			wait until rising_edge(clk);

			PA <= "11000010";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "01011000";
			PB <= "01000010";
			wait until rising_edge(clk);

			PA <= "01010011";
			PB <= "00001001";
			wait until rising_edge(clk);

			PA <= "00111110";
			PB <= "00100000";
			wait until rising_edge(clk);

			PA <= "10011010";
			PB <= "10010000";
			wait until rising_edge(clk);

			PA <= "10111000";
			PB <= "10100101";
			wait until rising_edge(clk);

			PA <= "00010100";
			PB <= "11010100";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "00011011";
			wait until rising_edge(clk);

			PA <= "11111110";
			PB <= "00111110";
			wait until rising_edge(clk);

			PA <= "11010111";
			PB <= "10011010";
			wait until rising_edge(clk);

			PA <= "00110111";
			PB <= "10001000";
			wait until rising_edge(clk);

			PA <= "01000110";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "00001000";
			PB <= "01000111";
			wait until rising_edge(clk);

			PA <= "01100101";
			PB <= "11011001";
			wait until rising_edge(clk);

			PA <= "00011110";
			PB <= "10001110";
			wait until rising_edge(clk);

			PA <= "10011110";
			PB <= "11000101";
			wait until rising_edge(clk);

			PA <= "11101100";
			PB <= "00010111";
			wait until rising_edge(clk);

			PA <= "00010010";
			PB <= "00110100";
			wait until rising_edge(clk);

			PA <= "11011010";
			PB <= "11000111";
			wait until rising_edge(clk);

			PA <= "00001100";
			PB <= "11010101";
			wait until rising_edge(clk);

			PA <= "11101011";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "00100111";
			PB <= "10011100";
			wait until rising_edge(clk);

			PA <= "11011111";
			PB <= "00000100";
			wait until rising_edge(clk);

			PA <= "01111111";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "00000111";
			PB <= "00100100";
			wait until rising_edge(clk);

			PA <= "01110011";
			PB <= "00111101";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "00101011";
			wait until rising_edge(clk);

			PA <= "01101110";
			PB <= "01010110";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "00101100";
			wait until rising_edge(clk);

			PA <= "11000111";
			PB <= "01001110";
			wait until rising_edge(clk);

			PA <= "01100011";
			PB <= "10011110";
			wait until rising_edge(clk);

			PA <= "11010000";
			PB <= "00001010";
			wait until rising_edge(clk);

			PA <= "00010100";
			PB <= "11011110";
			wait until rising_edge(clk);

			PA <= "00100000";
			PB <= "10000110";
			wait until rising_edge(clk);

			PA <= "11001111";
			PB <= "01011111";
			wait until rising_edge(clk);

			PA <= "01111000";
			PB <= "00011101";
			wait until rising_edge(clk);

			PA <= "11110101";
			PB <= "00010000";
			wait until rising_edge(clk);

			PA <= "00100101";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "11101001";
			PB <= "01001101";
			wait until rising_edge(clk);

			PA <= "10001101";
			PB <= "00000101";
			wait until rising_edge(clk);

			PA <= "11110001";
			PB <= "10100100";
			wait until rising_edge(clk);

			PA <= "10101001";
			PB <= "11110100";
			wait until rising_edge(clk);

			PA <= "10001000";
			PB <= "11001000";
			wait until rising_edge(clk);

			PA <= "00000001";
			PB <= "11111100";
			wait until rising_edge(clk);

			PA <= "11111100";
			PB <= "11110110";
			wait until rising_edge(clk);

			PA <= "01010111";
			PB <= "11001001";
			wait until rising_edge(clk);

			PA <= "10101101";
			PB <= "01110111";
			wait until rising_edge(clk);

			PA <= "10011110";
			PB <= "00011100";
			wait until rising_edge(clk);

			PA <= "11001010";
			PB <= "11111100";
			wait until rising_edge(clk);

			----------------------------------


	  		wait for 3330 ns;
	  		testing <= False;
	  		wait;
	  	end process;

	  	
	  	drive_rst: process
	  	begin
	  		reset <= '0';
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		reset <= '1';
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		reset <= '0';
	  		wait for 1500 ns;
	  		reset <= '1';
	  		wait for 330 ns;
	  		reset <= '0';
	  		wait for 2000 ns;
	  		reset <= '1';
	  		wait for 100 ns;
	  		reset <= '0';
	  		wait for 3000 ns;

	  		wait;
	  	end process;



	  	drive_en : process
	  	begin
	  		enable <= '1';
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		enable <= '0';
	  		wait until rising_edge(clk);
	  		wait until rising_edge(clk);
	  		enable <= '1';
	  		wait for 3000 ns;
	  		enable <= '0';
	  		wait for 200 ns;
	  		enable <= '1';
	  		wait for 2400 ns;
	  	end process;

end architecture;

